module kuznechik_cipher(
    input  logic         clk_i,     // Тактовый сигнал
    input  logic         resetn_i,  // Синхронный сигнал сброса с активным уровнем LOW
    input  logic         request_i, // Сигнал запроса на начало шифрования
    input  logic         ack_i,     // Сигнал подтверждения приема зашифрованных данных
    input  logic [127:0] data_i,    // Шифруемые данные

    output logic         busy_o,    // Сигнал, сообщающий о невозможности приёма
                                    // очередного запроса на шифрование, поскольку
                                    // модуль в процессе шифрования предыдущего
                                    // запроса
    output logic         valid_o,   // Сигнал готовности зашифрованных данных
    output logic [127:0] data_o     // Зашифрованные данные
);

  // Добавьте свой модуль сюда

endmodule
